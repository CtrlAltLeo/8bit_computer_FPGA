// Top level module with bus and submodules

module eightbit_computer(
	bus, // 8 bit wide bus
);

inout [7:0] bus;



endmodule
